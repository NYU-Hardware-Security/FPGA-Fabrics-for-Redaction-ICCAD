//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed May 26 01:10:41 2021
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
//`default_nettype none

// ----- Verilog module for fpga_top -----
module fpga_top(prog_clk,
                Test_en,
                IO_ISOL_N,
                clk,
                gfpga_pad_EMBEDDED_IO_HD_SOC_IN,
                gfpga_pad_EMBEDDED_IO_HD_SOC_OUT,
                gfpga_pad_EMBEDDED_IO_HD_SOC_DIR,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] Test_en;
//----- GLOBAL PORTS -----
input [0:0] IO_ISOL_N;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPIN PORTS -----
input [0:59] gfpga_pad_EMBEDDED_IO_HD_SOC_IN;
//----- GPOUT PORTS -----
output [0:59] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT;
//----- GPOUT PORTS -----
output [0:59] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:13] cbx_1__0__0_chanx_left_out;
wire [0:13] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:13] cbx_1__0__1_chanx_left_out;
wire [0:13] cbx_1__0__1_chanx_right_out;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__2_ccff_tail;
wire [0:13] cbx_1__0__2_chanx_left_out;
wire [0:13] cbx_1__0__2_chanx_right_out;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__3_ccff_tail;
wire [0:13] cbx_1__0__3_chanx_left_out;
wire [0:13] cbx_1__0__3_chanx_right_out;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__4_ccff_tail;
wire [0:13] cbx_1__0__4_chanx_left_out;
wire [0:13] cbx_1__0__4_chanx_right_out;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__0_ccff_tail;
wire [0:13] cbx_1__1__0_chanx_left_out;
wire [0:13] cbx_1__1__0_chanx_right_out;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__10_ccff_tail;
wire [0:13] cbx_1__1__10_chanx_left_out;
wire [0:13] cbx_1__1__10_chanx_right_out;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__11_ccff_tail;
wire [0:13] cbx_1__1__11_chanx_left_out;
wire [0:13] cbx_1__1__11_chanx_right_out;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__12_ccff_tail;
wire [0:13] cbx_1__1__12_chanx_left_out;
wire [0:13] cbx_1__1__12_chanx_right_out;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__13_ccff_tail;
wire [0:13] cbx_1__1__13_chanx_left_out;
wire [0:13] cbx_1__1__13_chanx_right_out;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__14_ccff_tail;
wire [0:13] cbx_1__1__14_chanx_left_out;
wire [0:13] cbx_1__1__14_chanx_right_out;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__15_ccff_tail;
wire [0:13] cbx_1__1__15_chanx_left_out;
wire [0:13] cbx_1__1__15_chanx_right_out;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__16_ccff_tail;
wire [0:13] cbx_1__1__16_chanx_left_out;
wire [0:13] cbx_1__1__16_chanx_right_out;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__17_ccff_tail;
wire [0:13] cbx_1__1__17_chanx_left_out;
wire [0:13] cbx_1__1__17_chanx_right_out;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__18_ccff_tail;
wire [0:13] cbx_1__1__18_chanx_left_out;
wire [0:13] cbx_1__1__18_chanx_right_out;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__19_ccff_tail;
wire [0:13] cbx_1__1__19_chanx_left_out;
wire [0:13] cbx_1__1__19_chanx_right_out;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__1_ccff_tail;
wire [0:13] cbx_1__1__1_chanx_left_out;
wire [0:13] cbx_1__1__1_chanx_right_out;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__2_ccff_tail;
wire [0:13] cbx_1__1__2_chanx_left_out;
wire [0:13] cbx_1__1__2_chanx_right_out;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__3_ccff_tail;
wire [0:13] cbx_1__1__3_chanx_left_out;
wire [0:13] cbx_1__1__3_chanx_right_out;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__4_ccff_tail;
wire [0:13] cbx_1__1__4_chanx_left_out;
wire [0:13] cbx_1__1__4_chanx_right_out;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__5_ccff_tail;
wire [0:13] cbx_1__1__5_chanx_left_out;
wire [0:13] cbx_1__1__5_chanx_right_out;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__6_ccff_tail;
wire [0:13] cbx_1__1__6_chanx_left_out;
wire [0:13] cbx_1__1__6_chanx_right_out;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__7_ccff_tail;
wire [0:13] cbx_1__1__7_chanx_left_out;
wire [0:13] cbx_1__1__7_chanx_right_out;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__8_ccff_tail;
wire [0:13] cbx_1__1__8_chanx_left_out;
wire [0:13] cbx_1__1__8_chanx_right_out;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__9_ccff_tail;
wire [0:13] cbx_1__1__9_chanx_left_out;
wire [0:13] cbx_1__1__9_chanx_right_out;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__5__0_ccff_tail;
wire [0:13] cbx_1__5__0_chanx_left_out;
wire [0:13] cbx_1__5__0_chanx_right_out;
wire [0:0] cbx_1__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__5__1_ccff_tail;
wire [0:13] cbx_1__5__1_chanx_left_out;
wire [0:13] cbx_1__5__1_chanx_right_out;
wire [0:0] cbx_1__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__5__2_ccff_tail;
wire [0:13] cbx_1__5__2_chanx_left_out;
wire [0:13] cbx_1__5__2_chanx_right_out;
wire [0:0] cbx_1__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__5__3_ccff_tail;
wire [0:13] cbx_1__5__3_chanx_left_out;
wire [0:13] cbx_1__5__3_chanx_right_out;
wire [0:0] cbx_1__5__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__5__4_ccff_tail;
wire [0:13] cbx_1__5__4_chanx_left_out;
wire [0:13] cbx_1__5__4_chanx_right_out;
wire [0:0] cbx_1__5__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:13] cby_0__1__0_chany_bottom_out;
wire [0:13] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:13] cby_0__1__1_chany_bottom_out;
wire [0:13] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__2_ccff_tail;
wire [0:13] cby_0__1__2_chany_bottom_out;
wire [0:13] cby_0__1__2_chany_top_out;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__3_ccff_tail;
wire [0:13] cby_0__1__3_chany_bottom_out;
wire [0:13] cby_0__1__3_chany_top_out;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__4_ccff_tail;
wire [0:13] cby_0__1__4_chany_bottom_out;
wire [0:13] cby_0__1__4_chany_top_out;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_1__1__0_ccff_tail;
wire [0:13] cby_1__1__0_chany_bottom_out;
wire [0:13] cby_1__1__0_chany_top_out;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__10_ccff_tail;
wire [0:13] cby_1__1__10_chany_bottom_out;
wire [0:13] cby_1__1__10_chany_top_out;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__11_ccff_tail;
wire [0:13] cby_1__1__11_chany_bottom_out;
wire [0:13] cby_1__1__11_chany_top_out;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__12_ccff_tail;
wire [0:13] cby_1__1__12_chany_bottom_out;
wire [0:13] cby_1__1__12_chany_top_out;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__13_ccff_tail;
wire [0:13] cby_1__1__13_chany_bottom_out;
wire [0:13] cby_1__1__13_chany_top_out;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__14_ccff_tail;
wire [0:13] cby_1__1__14_chany_bottom_out;
wire [0:13] cby_1__1__14_chany_top_out;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__15_ccff_tail;
wire [0:13] cby_1__1__15_chany_bottom_out;
wire [0:13] cby_1__1__15_chany_top_out;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__16_ccff_tail;
wire [0:13] cby_1__1__16_chany_bottom_out;
wire [0:13] cby_1__1__16_chany_top_out;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__17_ccff_tail;
wire [0:13] cby_1__1__17_chany_bottom_out;
wire [0:13] cby_1__1__17_chany_top_out;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__18_ccff_tail;
wire [0:13] cby_1__1__18_chany_bottom_out;
wire [0:13] cby_1__1__18_chany_top_out;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__19_ccff_tail;
wire [0:13] cby_1__1__19_chany_bottom_out;
wire [0:13] cby_1__1__19_chany_top_out;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__1_ccff_tail;
wire [0:13] cby_1__1__1_chany_bottom_out;
wire [0:13] cby_1__1__1_chany_top_out;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__2_ccff_tail;
wire [0:13] cby_1__1__2_chany_bottom_out;
wire [0:13] cby_1__1__2_chany_top_out;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__3_ccff_tail;
wire [0:13] cby_1__1__3_chany_bottom_out;
wire [0:13] cby_1__1__3_chany_top_out;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__4_ccff_tail;
wire [0:13] cby_1__1__4_chany_bottom_out;
wire [0:13] cby_1__1__4_chany_top_out;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__5_ccff_tail;
wire [0:13] cby_1__1__5_chany_bottom_out;
wire [0:13] cby_1__1__5_chany_top_out;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__6_ccff_tail;
wire [0:13] cby_1__1__6_chany_bottom_out;
wire [0:13] cby_1__1__6_chany_top_out;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__7_ccff_tail;
wire [0:13] cby_1__1__7_chany_bottom_out;
wire [0:13] cby_1__1__7_chany_top_out;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__8_ccff_tail;
wire [0:13] cby_1__1__8_chany_bottom_out;
wire [0:13] cby_1__1__8_chany_top_out;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__9_ccff_tail;
wire [0:13] cby_1__1__9_chany_bottom_out;
wire [0:13] cby_1__1__9_chany_top_out;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_5__1__0_ccff_tail;
wire [0:13] cby_5__1__0_chany_bottom_out;
wire [0:13] cby_5__1__0_chany_top_out;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_5__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_5__1__1_ccff_tail;
wire [0:13] cby_5__1__1_chany_bottom_out;
wire [0:13] cby_5__1__1_chany_top_out;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_5__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_5__1__2_ccff_tail;
wire [0:13] cby_5__1__2_chany_bottom_out;
wire [0:13] cby_5__1__2_chany_top_out;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_5__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_5__1__3_ccff_tail;
wire [0:13] cby_5__1__3_chany_bottom_out;
wire [0:13] cby_5__1__3_chany_top_out;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_5__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_5__1__4_ccff_tail;
wire [0:13] cby_5__1__4_chany_bottom_out;
wire [0:13] cby_5__1__4_chany_top_out;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_5__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] direct_interc_0_out;
wire [0:0] direct_interc_10_out;
wire [0:0] direct_interc_11_out;
wire [0:0] direct_interc_12_out;
wire [0:0] direct_interc_13_out;
wire [0:0] direct_interc_14_out;
wire [0:0] direct_interc_15_out;
wire [0:0] direct_interc_16_out;
wire [0:0] direct_interc_17_out;
wire [0:0] direct_interc_18_out;
wire [0:0] direct_interc_19_out;
wire [0:0] direct_interc_1_out;
wire [0:0] direct_interc_20_out;
wire [0:0] direct_interc_21_out;
wire [0:0] direct_interc_22_out;
wire [0:0] direct_interc_23_out;
wire [0:0] direct_interc_24_out;
wire [0:0] direct_interc_25_out;
wire [0:0] direct_interc_26_out;
wire [0:0] direct_interc_27_out;
wire [0:0] direct_interc_28_out;
wire [0:0] direct_interc_29_out;
wire [0:0] direct_interc_2_out;
wire [0:0] direct_interc_30_out;
wire [0:0] direct_interc_31_out;
wire [0:0] direct_interc_32_out;
wire [0:0] direct_interc_33_out;
wire [0:0] direct_interc_34_out;
wire [0:0] direct_interc_35_out;
wire [0:0] direct_interc_36_out;
wire [0:0] direct_interc_37_out;
wire [0:0] direct_interc_38_out;
wire [0:0] direct_interc_39_out;
wire [0:0] direct_interc_3_out;
wire [0:0] direct_interc_40_out;
wire [0:0] direct_interc_41_out;
wire [0:0] direct_interc_42_out;
wire [0:0] direct_interc_43_out;
wire [0:0] direct_interc_4_out;
wire [0:0] direct_interc_5_out;
wire [0:0] direct_interc_6_out;
wire [0:0] direct_interc_7_out;
wire [0:0] direct_interc_8_out;
wire [0:0] direct_interc_9_out;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_10_ccff_tail;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_11_ccff_tail;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_12_ccff_tail;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_13_ccff_tail;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_14_ccff_tail;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_15_ccff_tail;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_16_ccff_tail;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_17_ccff_tail;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_18_ccff_tail;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_19_ccff_tail;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_1__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
wire [0:0] grid_clb_1__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_1_ccff_tail;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_20_ccff_tail;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_21_ccff_tail;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_22_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_22_ccff_tail;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_23_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_23_ccff_tail;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_24_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_2__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_3__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_3_ccff_tail;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_4__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_4_ccff_tail;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_5__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_5_ccff_tail;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_6_ccff_tail;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_7_ccff_tail;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_8_ccff_tail;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_9_ccff_tail;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_io_bottom_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_2_ccff_tail;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_3_ccff_tail;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_4_ccff_tail;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_;
wire [0:0] grid_io_left_left_0_ccff_tail;
wire [0:0] grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_left_1_ccff_tail;
wire [0:0] grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_left_2_ccff_tail;
wire [0:0] grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_left_3_ccff_tail;
wire [0:0] grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_left_4_ccff_tail;
wire [0:0] grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_right_0_ccff_tail;
wire [0:0] grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_right_1_ccff_tail;
wire [0:0] grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_right_2_ccff_tail;
wire [0:0] grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_right_3_ccff_tail;
wire [0:0] grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_right_4_ccff_tail;
wire [0:0] grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_top_0_ccff_tail;
wire [0:0] grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_top_1_ccff_tail;
wire [0:0] grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_top_2_ccff_tail;
wire [0:0] grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_top_3_ccff_tail;
wire [0:0] grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_top_4_ccff_tail;
wire [0:0] sb_0__0__0_ccff_tail;
wire [0:13] sb_0__0__0_chanx_right_out;
wire [0:13] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:13] sb_0__1__0_chanx_right_out;
wire [0:13] sb_0__1__0_chany_bottom_out;
wire [0:13] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__1__1_ccff_tail;
wire [0:13] sb_0__1__1_chanx_right_out;
wire [0:13] sb_0__1__1_chany_bottom_out;
wire [0:13] sb_0__1__1_chany_top_out;
wire [0:0] sb_0__1__2_ccff_tail;
wire [0:13] sb_0__1__2_chanx_right_out;
wire [0:13] sb_0__1__2_chany_bottom_out;
wire [0:13] sb_0__1__2_chany_top_out;
wire [0:0] sb_0__1__3_ccff_tail;
wire [0:13] sb_0__1__3_chanx_right_out;
wire [0:13] sb_0__1__3_chany_bottom_out;
wire [0:13] sb_0__1__3_chany_top_out;
wire [0:0] sb_0__5__0_ccff_tail;
wire [0:13] sb_0__5__0_chanx_right_out;
wire [0:13] sb_0__5__0_chany_bottom_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:13] sb_1__0__0_chanx_left_out;
wire [0:13] sb_1__0__0_chanx_right_out;
wire [0:13] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__0__1_ccff_tail;
wire [0:13] sb_1__0__1_chanx_left_out;
wire [0:13] sb_1__0__1_chanx_right_out;
wire [0:13] sb_1__0__1_chany_top_out;
wire [0:0] sb_1__0__2_ccff_tail;
wire [0:13] sb_1__0__2_chanx_left_out;
wire [0:13] sb_1__0__2_chanx_right_out;
wire [0:13] sb_1__0__2_chany_top_out;
wire [0:0] sb_1__0__3_ccff_tail;
wire [0:13] sb_1__0__3_chanx_left_out;
wire [0:13] sb_1__0__3_chanx_right_out;
wire [0:13] sb_1__0__3_chany_top_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:13] sb_1__1__0_chanx_left_out;
wire [0:13] sb_1__1__0_chanx_right_out;
wire [0:13] sb_1__1__0_chany_bottom_out;
wire [0:13] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__1__10_ccff_tail;
wire [0:13] sb_1__1__10_chanx_left_out;
wire [0:13] sb_1__1__10_chanx_right_out;
wire [0:13] sb_1__1__10_chany_bottom_out;
wire [0:13] sb_1__1__10_chany_top_out;
wire [0:0] sb_1__1__11_ccff_tail;
wire [0:13] sb_1__1__11_chanx_left_out;
wire [0:13] sb_1__1__11_chanx_right_out;
wire [0:13] sb_1__1__11_chany_bottom_out;
wire [0:13] sb_1__1__11_chany_top_out;
wire [0:0] sb_1__1__12_ccff_tail;
wire [0:13] sb_1__1__12_chanx_left_out;
wire [0:13] sb_1__1__12_chanx_right_out;
wire [0:13] sb_1__1__12_chany_bottom_out;
wire [0:13] sb_1__1__12_chany_top_out;
wire [0:0] sb_1__1__13_ccff_tail;
wire [0:13] sb_1__1__13_chanx_left_out;
wire [0:13] sb_1__1__13_chanx_right_out;
wire [0:13] sb_1__1__13_chany_bottom_out;
wire [0:13] sb_1__1__13_chany_top_out;
wire [0:0] sb_1__1__14_ccff_tail;
wire [0:13] sb_1__1__14_chanx_left_out;
wire [0:13] sb_1__1__14_chanx_right_out;
wire [0:13] sb_1__1__14_chany_bottom_out;
wire [0:13] sb_1__1__14_chany_top_out;
wire [0:0] sb_1__1__15_ccff_tail;
wire [0:13] sb_1__1__15_chanx_left_out;
wire [0:13] sb_1__1__15_chanx_right_out;
wire [0:13] sb_1__1__15_chany_bottom_out;
wire [0:13] sb_1__1__15_chany_top_out;
wire [0:0] sb_1__1__1_ccff_tail;
wire [0:13] sb_1__1__1_chanx_left_out;
wire [0:13] sb_1__1__1_chanx_right_out;
wire [0:13] sb_1__1__1_chany_bottom_out;
wire [0:13] sb_1__1__1_chany_top_out;
wire [0:0] sb_1__1__2_ccff_tail;
wire [0:13] sb_1__1__2_chanx_left_out;
wire [0:13] sb_1__1__2_chanx_right_out;
wire [0:13] sb_1__1__2_chany_bottom_out;
wire [0:13] sb_1__1__2_chany_top_out;
wire [0:0] sb_1__1__3_ccff_tail;
wire [0:13] sb_1__1__3_chanx_left_out;
wire [0:13] sb_1__1__3_chanx_right_out;
wire [0:13] sb_1__1__3_chany_bottom_out;
wire [0:13] sb_1__1__3_chany_top_out;
wire [0:0] sb_1__1__4_ccff_tail;
wire [0:13] sb_1__1__4_chanx_left_out;
wire [0:13] sb_1__1__4_chanx_right_out;
wire [0:13] sb_1__1__4_chany_bottom_out;
wire [0:13] sb_1__1__4_chany_top_out;
wire [0:0] sb_1__1__5_ccff_tail;
wire [0:13] sb_1__1__5_chanx_left_out;
wire [0:13] sb_1__1__5_chanx_right_out;
wire [0:13] sb_1__1__5_chany_bottom_out;
wire [0:13] sb_1__1__5_chany_top_out;
wire [0:0] sb_1__1__6_ccff_tail;
wire [0:13] sb_1__1__6_chanx_left_out;
wire [0:13] sb_1__1__6_chanx_right_out;
wire [0:13] sb_1__1__6_chany_bottom_out;
wire [0:13] sb_1__1__6_chany_top_out;
wire [0:0] sb_1__1__7_ccff_tail;
wire [0:13] sb_1__1__7_chanx_left_out;
wire [0:13] sb_1__1__7_chanx_right_out;
wire [0:13] sb_1__1__7_chany_bottom_out;
wire [0:13] sb_1__1__7_chany_top_out;
wire [0:0] sb_1__1__8_ccff_tail;
wire [0:13] sb_1__1__8_chanx_left_out;
wire [0:13] sb_1__1__8_chanx_right_out;
wire [0:13] sb_1__1__8_chany_bottom_out;
wire [0:13] sb_1__1__8_chany_top_out;
wire [0:0] sb_1__1__9_ccff_tail;
wire [0:13] sb_1__1__9_chanx_left_out;
wire [0:13] sb_1__1__9_chanx_right_out;
wire [0:13] sb_1__1__9_chany_bottom_out;
wire [0:13] sb_1__1__9_chany_top_out;
wire [0:0] sb_1__5__0_ccff_tail;
wire [0:13] sb_1__5__0_chanx_left_out;
wire [0:13] sb_1__5__0_chanx_right_out;
wire [0:13] sb_1__5__0_chany_bottom_out;
wire [0:0] sb_1__5__1_ccff_tail;
wire [0:13] sb_1__5__1_chanx_left_out;
wire [0:13] sb_1__5__1_chanx_right_out;
wire [0:13] sb_1__5__1_chany_bottom_out;
wire [0:0] sb_1__5__2_ccff_tail;
wire [0:13] sb_1__5__2_chanx_left_out;
wire [0:13] sb_1__5__2_chanx_right_out;
wire [0:13] sb_1__5__2_chany_bottom_out;
wire [0:0] sb_1__5__3_ccff_tail;
wire [0:13] sb_1__5__3_chanx_left_out;
wire [0:13] sb_1__5__3_chanx_right_out;
wire [0:13] sb_1__5__3_chany_bottom_out;
wire [0:0] sb_5__0__0_ccff_tail;
wire [0:13] sb_5__0__0_chanx_left_out;
wire [0:13] sb_5__0__0_chany_top_out;
wire [0:0] sb_5__1__0_ccff_tail;
wire [0:13] sb_5__1__0_chanx_left_out;
wire [0:13] sb_5__1__0_chany_bottom_out;
wire [0:13] sb_5__1__0_chany_top_out;
wire [0:0] sb_5__1__1_ccff_tail;
wire [0:13] sb_5__1__1_chanx_left_out;
wire [0:13] sb_5__1__1_chany_bottom_out;
wire [0:13] sb_5__1__1_chany_top_out;
wire [0:0] sb_5__1__2_ccff_tail;
wire [0:13] sb_5__1__2_chanx_left_out;
wire [0:13] sb_5__1__2_chany_bottom_out;
wire [0:13] sb_5__1__2_chany_top_out;
wire [0:0] sb_5__1__3_ccff_tail;
wire [0:13] sb_5__1__3_chanx_left_out;
wire [0:13] sb_5__1__3_chany_bottom_out;
wire [0:13] sb_5__1__3_chany_top_out;
wire [0:0] sb_5__5__0_ccff_tail;
wire [0:13] sb_5__5__0_chanx_left_out;
wire [0:13] sb_5__5__0_chany_bottom_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_clb grid_clb_1__1_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_0_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_20_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__2_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_1_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_21_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_1__3_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_2_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_22_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_1__4_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_3_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_23_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_3_ccff_tail));

	grid_clb grid_clb_1__5_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_1__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_2__1_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_4_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_24_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_2__2_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_5_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_25_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_2__3_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_6_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_26_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_7_ccff_tail));

	grid_clb grid_clb_2__4_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_7_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_27_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_8_ccff_tail));

	grid_clb grid_clb_2__5_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_2__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_40_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_9_ccff_tail));

	grid_clb grid_clb_3__1_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_8_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_28_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_10_ccff_tail));

	grid_clb grid_clb_3__2_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_9_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_29_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_11_ccff_tail));

	grid_clb grid_clb_3__3_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_10_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_30_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_12_ccff_tail));

	grid_clb grid_clb_3__4_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_11_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_31_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_13_ccff_tail));

	grid_clb grid_clb_3__5_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_3__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_41_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_14_ccff_tail));

	grid_clb grid_clb_4__1_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_12_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_32_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_15_ccff_tail));

	grid_clb grid_clb_4__2_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_13_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_33_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_16_ccff_tail));

	grid_clb grid_clb_4__3_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_14_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_34_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_17_ccff_tail));

	grid_clb grid_clb_4__4_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_15_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_35_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__18_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_18_ccff_tail));

	grid_clb grid_clb_4__5_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_4__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_42_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__19_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_19_ccff_tail));

	grid_clb grid_clb_5__1_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_16_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_36_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_5__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_20_ccff_tail));

	grid_clb grid_clb_5__2_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_17_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_37_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_5__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_21_ccff_tail));

	grid_clb grid_clb_5__3_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_18_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_38_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_5__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_22_ccff_tail));

	grid_clb grid_clb_5__4_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_19_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_39_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_5__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_23_ccff_tail));

	grid_clb grid_clb_5__5_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_5__5__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_43_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_5__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(ccff_tail));

	grid_io_top_top grid_io_top_top_1__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__5__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_0_ccff_tail));

	grid_io_top_top grid_io_top_top_2__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__5__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_1_ccff_tail));

	grid_io_top_top grid_io_top_top_3__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__5__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_2_ccff_tail));

	grid_io_top_top grid_io_top_top_4__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__5__3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_3_ccff_tail));

	grid_io_top_top grid_io_top_top_5__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__5__4_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_4_ccff_tail));

	grid_io_right_right grid_io_right_right_6__5_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_0_ccff_tail));

	grid_io_right_right grid_io_right_right_6__4_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_1_ccff_tail));

	grid_io_right_right grid_io_right_right_6__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_2_ccff_tail));

	grid_io_right_right grid_io_right_right_6__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_4_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_3_ccff_tail));

	grid_io_right_right grid_io_right_right_6__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_4_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_5__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10:18]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10:18]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10:18]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_0_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_4__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19:27]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19:27]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19:27]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_1_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_3__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28:36]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28:36]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28:36]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_2_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_2__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37:45]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37:45]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37:45]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_3_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_1__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46:54]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46:54]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46:54]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_4_ccff_tail));

	grid_io_left_left grid_io_left_left_0__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_0_ccff_tail));

	grid_io_left_left grid_io_left_left_0__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_1_ccff_tail));

	grid_io_left_left grid_io_left_left_0__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_2_ccff_tail));

	grid_io_left_left grid_io_left_left_0__4_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_3_ccff_tail));

	grid_io_left_left grid_io_left_left_0__5_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__4_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_4_ccff_tail));

	sb_0__0_ sb_0__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_head(grid_io_left_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:13]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:13]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_left_2_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:13]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:13]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:13]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__1_ sb_0__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_left_3_ccff_tail),
		.chany_top_out(sb_0__1__1_chany_top_out[0:13]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:13]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:13]),
		.ccff_tail(sb_0__1__1_ccff_tail));

	sb_0__1_ sb_0__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_left_4_ccff_tail),
		.chany_top_out(sb_0__1__2_chany_top_out[0:13]),
		.chanx_right_out(sb_0__1__2_chanx_right_out[0:13]),
		.chany_bottom_out(sb_0__1__2_chany_bottom_out[0:13]),
		.ccff_tail(sb_0__1__2_ccff_tail));

	sb_0__1_ sb_0__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__4_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(sb_0__5__0_ccff_tail),
		.chany_top_out(sb_0__1__3_chany_top_out[0:13]),
		.chanx_right_out(sb_0__1__3_chanx_right_out[0:13]),
		.chany_bottom_out(sb_0__1__3_chany_bottom_out[0:13]),
		.ccff_tail(sb_0__1__3_ccff_tail));

	sb_0__5_ sb_0__5_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__5__0_chanx_left_out[0:13]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_top_top_0_ccff_tail),
		.chanx_right_out(sb_0__5__0_chanx_right_out[0:13]),
		.chany_bottom_out(sb_0__5__0_chany_bottom_out[0:13]),
		.ccff_tail(sb_0__5__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_head(grid_io_left_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:13]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:13]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:13]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:13]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:13]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:13]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__0_ sb_3__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__10_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_1__0__2_chany_top_out[0:13]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:13]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:13]),
		.ccff_tail(sb_1__0__2_ccff_tail));

	sb_1__0_ sb_4__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__15_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_head(grid_clb_10_ccff_tail),
		.chany_top_out(sb_1__0__3_chany_top_out[0:13]),
		.chanx_right_out(sb_1__0__3_chanx_right_out[0:13]),
		.chanx_left_out(sb_1__0__3_chanx_left_out[0:13]),
		.ccff_tail(sb_1__0__3_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__4_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_1__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__5_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__1_ sb_1__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__6_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_8_ccff_tail),
		.chany_top_out(sb_1__1__2_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__2_ccff_tail));

	sb_1__1_ sb_1__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__7_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_3_ccff_tail),
		.chany_top_out(sb_1__1__3_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__3_ccff_tail));

	sb_1__1_ sb_2__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__8_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__4_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_11_ccff_tail),
		.chany_top_out(sb_1__1__4_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__4_ccff_tail));

	sb_1__1_ sb_2__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__9_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__5_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__1__5_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__5_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__5_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__5_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__5_ccff_tail));

	sb_1__1_ sb_2__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__8_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__10_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__6_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_13_ccff_tail),
		.chany_top_out(sb_1__1__6_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__6_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__6_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__6_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__6_ccff_tail));

	sb_1__1_ sb_2__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__9_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__11_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__7_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__1__7_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__7_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__7_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__7_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__7_ccff_tail));

	sb_1__1_ sb_3__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__11_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__12_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__8_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_16_ccff_tail),
		.chany_top_out(sb_1__1__8_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__8_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__8_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__8_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__8_ccff_tail));

	sb_1__1_ sb_3__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__12_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__13_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__9_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_7_ccff_tail),
		.chany_top_out(sb_1__1__9_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__9_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__9_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__9_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__9_ccff_tail));

	sb_1__1_ sb_3__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__13_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__14_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__12_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__10_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_18_ccff_tail),
		.chany_top_out(sb_1__1__10_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__10_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__10_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__10_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__10_ccff_tail));

	sb_1__1_ sb_3__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__14_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__15_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__13_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__11_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_9_ccff_tail),
		.chany_top_out(sb_1__1__11_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__11_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__11_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__11_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__11_ccff_tail));

	sb_1__1_ sb_4__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__16_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__16_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__15_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__12_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_21_ccff_tail),
		.chany_top_out(sb_1__1__12_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__12_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__12_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__12_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__12_ccff_tail));

	sb_1__1_ sb_4__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__17_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__17_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__16_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__13_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_12_ccff_tail),
		.chany_top_out(sb_1__1__13_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__13_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__13_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__13_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__13_ccff_tail));

	sb_1__1_ sb_4__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__18_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__18_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__17_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__14_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_23_ccff_tail),
		.chany_top_out(sb_1__1__14_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__14_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__14_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__14_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__14_ccff_tail));

	sb_1__1_ sb_4__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__19_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__19_chanx_left_out[0:13]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__18_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__15_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_14_ccff_tail),
		.chany_top_out(sb_1__1__15_chany_top_out[0:13]),
		.chanx_right_out(sb_1__1__15_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__1__15_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__1__15_chanx_left_out[0:13]),
		.ccff_tail(sb_1__1__15_ccff_tail));

	sb_1__5_ sb_1__5_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__5__1_chanx_left_out[0:13]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__5__0_chanx_right_out[0:13]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_1_ccff_tail),
		.chanx_right_out(sb_1__5__0_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__5__0_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__5__0_chanx_left_out[0:13]),
		.ccff_tail(sb_1__5__0_ccff_tail));

	sb_1__5_ sb_2__5_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__5__2_chanx_left_out[0:13]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__5__1_chanx_right_out[0:13]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_2_ccff_tail),
		.chanx_right_out(sb_1__5__1_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__5__1_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__5__1_chanx_left_out[0:13]),
		.ccff_tail(sb_1__5__1_ccff_tail));

	sb_1__5_ sb_3__5_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__5__3_chanx_left_out[0:13]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__14_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__5__2_chanx_right_out[0:13]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_3_ccff_tail),
		.chanx_right_out(sb_1__5__2_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__5__2_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__5__2_chanx_left_out[0:13]),
		.ccff_tail(sb_1__5__2_ccff_tail));

	sb_1__5_ sb_4__5_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__5__4_chanx_left_out[0:13]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__19_chany_top_out[0:13]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__5__3_chanx_right_out[0:13]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_4_ccff_tail),
		.chanx_right_out(sb_1__5__3_chanx_right_out[0:13]),
		.chany_bottom_out(sb_1__5__3_chany_bottom_out[0:13]),
		.chanx_left_out(sb_1__5__3_chanx_left_out[0:13]),
		.ccff_tail(sb_1__5__3_ccff_tail));

	sb_5__0_ sb_5__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_5__1__0_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_),
		.ccff_head(grid_clb_15_ccff_tail),
		.chany_top_out(sb_5__0__0_chany_top_out[0:13]),
		.chanx_left_out(sb_5__0__0_chanx_left_out[0:13]),
		.ccff_tail(sb_5__0__0_ccff_tail));

	sb_5__1_ sb_5__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_5__1__1_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_5__1__0_chany_top_out[0:13]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__16_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_20_ccff_tail),
		.chany_top_out(sb_5__1__0_chany_top_out[0:13]),
		.chany_bottom_out(sb_5__1__0_chany_bottom_out[0:13]),
		.chanx_left_out(sb_5__1__0_chanx_left_out[0:13]),
		.ccff_tail(sb_5__1__0_ccff_tail));

	sb_5__1_ sb_5__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_5__1__2_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_5__1__1_chany_top_out[0:13]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__17_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_17_ccff_tail),
		.chany_top_out(sb_5__1__1_chany_top_out[0:13]),
		.chany_bottom_out(sb_5__1__1_chany_bottom_out[0:13]),
		.chanx_left_out(sb_5__1__1_chanx_left_out[0:13]),
		.ccff_tail(sb_5__1__1_ccff_tail));

	sb_5__1_ sb_5__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_5__1__3_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_5__1__2_chany_top_out[0:13]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__18_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_22_ccff_tail),
		.chany_top_out(sb_5__1__2_chany_top_out[0:13]),
		.chany_bottom_out(sb_5__1__2_chany_bottom_out[0:13]),
		.chanx_left_out(sb_5__1__2_chanx_left_out[0:13]),
		.ccff_tail(sb_5__1__2_ccff_tail));

	sb_5__1_ sb_5__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_5__1__4_chany_bottom_out[0:13]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_5__1__3_chany_top_out[0:13]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__19_chanx_right_out[0:13]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_19_ccff_tail),
		.chany_top_out(sb_5__1__3_chany_top_out[0:13]),
		.chany_bottom_out(sb_5__1__3_chany_bottom_out[0:13]),
		.chanx_left_out(sb_5__1__3_chanx_left_out[0:13]),
		.ccff_tail(sb_5__1__3_ccff_tail));

	sb_5__5_ sb_5__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_5__1__4_chany_top_out[0:13]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__5__4_chanx_right_out[0:13]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_right_right_0_ccff_tail),
		.chany_bottom_out(sb_5__5__0_chany_bottom_out[0:13]),
		.chanx_left_out(sb_5__5__0_chanx_left_out[0:13]),
		.ccff_tail(sb_5__5__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:13]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:13]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:13]),
		.ccff_head(sb_1__0__2_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__0_ cbx_4__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__0__3_chanx_left_out[0:13]),
		.ccff_head(sb_1__0__3_ccff_tail),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__3_ccff_tail));

	cbx_1__0_ cbx_5__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__3_chanx_right_out[0:13]),
		.chanx_right_in(sb_5__0__0_chanx_left_out[0:13]),
		.ccff_head(sb_5__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__4_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__0_ccff_tail));

	cbx_1__1_ cbx_1__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__1_ccff_tail));

	cbx_1__1_ cbx_1__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__2_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__2_ccff_tail));

	cbx_1__1_ cbx_1__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__3_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__3_ccff_tail),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__3_ccff_tail));

	cbx_1__1_ cbx_2__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__4_ccff_tail),
		.chanx_left_out(cbx_1__1__4_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__4_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__4_ccff_tail));

	cbx_1__1_ cbx_2__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__5_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__5_ccff_tail),
		.chanx_left_out(cbx_1__1__5_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__5_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__5_ccff_tail));

	cbx_1__1_ cbx_2__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__6_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__6_ccff_tail),
		.chanx_left_out(cbx_1__1__6_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__6_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__6_ccff_tail));

	cbx_1__1_ cbx_2__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__7_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__7_ccff_tail),
		.chanx_left_out(cbx_1__1__7_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__7_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__7_ccff_tail));

	cbx_1__1_ cbx_3__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__4_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__8_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__8_ccff_tail),
		.chanx_left_out(cbx_1__1__8_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__8_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__8_ccff_tail));

	cbx_1__1_ cbx_3__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__5_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__9_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__9_ccff_tail),
		.chanx_left_out(cbx_1__1__9_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__9_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__9_ccff_tail));

	cbx_1__1_ cbx_3__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__6_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__10_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__10_ccff_tail),
		.chanx_left_out(cbx_1__1__10_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__10_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__10_ccff_tail));

	cbx_1__1_ cbx_3__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__7_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__11_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__11_ccff_tail),
		.chanx_left_out(cbx_1__1__11_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__11_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__11_ccff_tail));

	cbx_1__1_ cbx_4__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__8_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__12_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__12_ccff_tail),
		.chanx_left_out(cbx_1__1__12_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__12_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__12_ccff_tail));

	cbx_1__1_ cbx_4__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__9_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__13_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__13_ccff_tail),
		.chanx_left_out(cbx_1__1__13_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__13_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__13_ccff_tail));

	cbx_1__1_ cbx_4__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__10_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__14_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__14_ccff_tail),
		.chanx_left_out(cbx_1__1__14_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__14_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__14_ccff_tail));

	cbx_1__1_ cbx_4__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__11_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__1__15_chanx_left_out[0:13]),
		.ccff_head(sb_1__1__15_ccff_tail),
		.chanx_left_out(cbx_1__1__15_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__15_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__15_ccff_tail));

	cbx_1__1_ cbx_5__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__12_chanx_right_out[0:13]),
		.chanx_right_in(sb_5__1__0_chanx_left_out[0:13]),
		.ccff_head(sb_5__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__16_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__16_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__16_ccff_tail));

	cbx_1__1_ cbx_5__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__13_chanx_right_out[0:13]),
		.chanx_right_in(sb_5__1__1_chanx_left_out[0:13]),
		.ccff_head(sb_5__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__17_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__17_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__17_ccff_tail));

	cbx_1__1_ cbx_5__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__14_chanx_right_out[0:13]),
		.chanx_right_in(sb_5__1__2_chanx_left_out[0:13]),
		.ccff_head(sb_5__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__18_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__18_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__18_ccff_tail));

	cbx_1__1_ cbx_5__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__15_chanx_right_out[0:13]),
		.chanx_right_in(sb_5__1__3_chanx_left_out[0:13]),
		.ccff_head(sb_5__1__3_ccff_tail),
		.chanx_left_out(cbx_1__1__19_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__1__19_chanx_right_out[0:13]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__19_ccff_tail));

	cbx_1__5_ cbx_1__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__5__0_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__5__0_chanx_left_out[0:13]),
		.ccff_head(sb_1__5__0_ccff_tail),
		.chanx_left_out(cbx_1__5__0_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__5__0_chanx_right_out[0:13]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__5__0_ccff_tail));

	cbx_1__5_ cbx_2__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__0_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__5__1_chanx_left_out[0:13]),
		.ccff_head(sb_1__5__1_ccff_tail),
		.chanx_left_out(cbx_1__5__1_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__5__1_chanx_right_out[0:13]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__5__1_ccff_tail));

	cbx_1__5_ cbx_3__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__1_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__5__2_chanx_left_out[0:13]),
		.ccff_head(sb_1__5__2_ccff_tail),
		.chanx_left_out(cbx_1__5__2_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__5__2_chanx_right_out[0:13]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__5__2_ccff_tail));

	cbx_1__5_ cbx_4__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__2_chanx_right_out[0:13]),
		.chanx_right_in(sb_1__5__3_chanx_left_out[0:13]),
		.ccff_head(sb_1__5__3_ccff_tail),
		.chanx_left_out(cbx_1__5__3_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__5__3_chanx_right_out[0:13]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__5__3_ccff_tail));

	cbx_1__5_ cbx_5__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__3_chanx_right_out[0:13]),
		.chanx_right_in(sb_5__5__0_chanx_left_out[0:13]),
		.ccff_head(sb_5__5__0_ccff_tail),
		.chanx_left_out(cbx_1__5__4_chanx_left_out[0:13]),
		.chanx_right_out(cbx_1__5__4_chanx_right_out[0:13]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__5__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__5__4_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:13]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:13]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:13]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:13]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:13]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:13]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_0__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:13]),
		.chany_top_in(sb_0__1__2_chany_bottom_out[0:13]),
		.ccff_head(sb_0__1__1_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:13]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_0__1_ cby_0__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__2_chany_top_out[0:13]),
		.chany_top_in(sb_0__1__3_chany_bottom_out[0:13]),
		.ccff_head(sb_0__1__2_ccff_tail),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:13]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__3_ccff_tail));

	cby_0__1_ cby_0__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__3_chany_top_out[0:13]),
		.chany_top_in(sb_0__5__0_chany_bottom_out[0:13]),
		.ccff_head(sb_0__1__3_ccff_tail),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:13]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__4_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__1_ cby_1__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__0_ccff_tail),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__1_ccff_tail));

	cby_1__1_ cby_1__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__1_ccff_tail),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__2_ccff_tail));

	cby_1__1_ cby_1__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__2_ccff_tail),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__3_ccff_tail));

	cby_1__1_ cby_1__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:13]),
		.chany_top_in(sb_1__5__0_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__3_ccff_tail),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__4_ccff_tail));

	cby_1__1_ cby_2__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__5_ccff_tail));

	cby_1__1_ cby_2__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__4_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__5_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__4_ccff_tail),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__6_ccff_tail));

	cby_1__1_ cby_2__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__5_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__6_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__5_ccff_tail),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__7_ccff_tail));

	cby_1__1_ cby_2__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__6_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__7_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__6_ccff_tail),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__8_ccff_tail));

	cby_1__1_ cby_2__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__7_chany_top_out[0:13]),
		.chany_top_in(sb_1__5__1_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__7_ccff_tail),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__9_ccff_tail));

	cby_1__1_ cby_3__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__8_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__10_ccff_tail));

	cby_1__1_ cby_3__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__8_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__9_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__8_ccff_tail),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__11_ccff_tail));

	cby_1__1_ cby_3__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__9_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__10_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__9_ccff_tail),
		.chany_bottom_out(cby_1__1__12_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__12_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__12_ccff_tail));

	cby_1__1_ cby_3__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__10_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__11_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__10_ccff_tail),
		.chany_bottom_out(cby_1__1__13_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__13_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__13_ccff_tail));

	cby_1__1_ cby_3__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__11_chany_top_out[0:13]),
		.chany_top_in(sb_1__5__2_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__11_ccff_tail),
		.chany_bottom_out(cby_1__1__14_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__14_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__14_ccff_tail));

	cby_1__1_ cby_4__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__3_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__12_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__0__3_ccff_tail),
		.chany_bottom_out(cby_1__1__15_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__15_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__15_ccff_tail));

	cby_1__1_ cby_4__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__12_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__13_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__12_ccff_tail),
		.chany_bottom_out(cby_1__1__16_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__16_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__16_ccff_tail));

	cby_1__1_ cby_4__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__13_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__14_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__13_ccff_tail),
		.chany_bottom_out(cby_1__1__17_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__17_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__17_ccff_tail));

	cby_1__1_ cby_4__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__14_chany_top_out[0:13]),
		.chany_top_in(sb_1__1__15_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__14_ccff_tail),
		.chany_bottom_out(cby_1__1__18_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__18_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__18_ccff_tail));

	cby_1__1_ cby_4__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__15_chany_top_out[0:13]),
		.chany_top_in(sb_1__5__3_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__15_ccff_tail),
		.chany_bottom_out(cby_1__1__19_chany_bottom_out[0:13]),
		.chany_top_out(cby_1__1__19_chany_top_out[0:13]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__19_ccff_tail));

	cby_5__1_ cby_5__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_5__0__0_chany_top_out[0:13]),
		.chany_top_in(sb_5__1__0_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__0__4_ccff_tail),
		.chany_bottom_out(cby_5__1__0_chany_bottom_out[0:13]),
		.chany_top_out(cby_5__1__0_chany_top_out[0:13]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_5__1__0_ccff_tail));

	cby_5__1_ cby_5__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_5__1__0_chany_top_out[0:13]),
		.chany_top_in(sb_5__1__1_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__16_ccff_tail),
		.chany_bottom_out(cby_5__1__1_chany_bottom_out[0:13]),
		.chany_top_out(cby_5__1__1_chany_top_out[0:13]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_5__1__1_ccff_tail));

	cby_5__1_ cby_5__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_5__1__1_chany_top_out[0:13]),
		.chany_top_in(sb_5__1__2_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__17_ccff_tail),
		.chany_bottom_out(cby_5__1__2_chany_bottom_out[0:13]),
		.chany_top_out(cby_5__1__2_chany_top_out[0:13]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_5__1__2_ccff_tail));

	cby_5__1_ cby_5__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_5__1__2_chany_top_out[0:13]),
		.chany_top_in(sb_5__1__3_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__18_ccff_tail),
		.chany_bottom_out(cby_5__1__3_chany_bottom_out[0:13]),
		.chany_top_out(cby_5__1__3_chany_top_out[0:13]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_5__1__3_ccff_tail));

	cby_5__1_ cby_5__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_5__1__3_chany_top_out[0:13]),
		.chany_top_in(sb_5__5__0_chany_bottom_out[0:13]),
		.ccff_head(cbx_1__1__19_ccff_tail),
		.chany_bottom_out(cby_5__1__4_chany_bottom_out[0:13]),
		.chany_top_out(cby_5__1__4_chany_top_out[0:13]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_5__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_5__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_5__1__4_ccff_tail));

	direct_interc direct_interc_0_ (
		.in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_0_out));

	direct_interc direct_interc_1_ (
		.in(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_1_out));

	direct_interc direct_interc_2_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_2_out));

	direct_interc direct_interc_3_ (
		.in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_3_out));

	direct_interc direct_interc_4_ (
		.in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_4_out));

	direct_interc direct_interc_5_ (
		.in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_5_out));

	direct_interc direct_interc_6_ (
		.in(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_6_out));

	direct_interc direct_interc_7_ (
		.in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_7_out));

	direct_interc direct_interc_8_ (
		.in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_8_out));

	direct_interc direct_interc_9_ (
		.in(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_9_out));

	direct_interc direct_interc_10_ (
		.in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_10_out));

	direct_interc direct_interc_11_ (
		.in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_11_out));

	direct_interc direct_interc_12_ (
		.in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_12_out));

	direct_interc direct_interc_13_ (
		.in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_13_out));

	direct_interc direct_interc_14_ (
		.in(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_14_out));

	direct_interc direct_interc_15_ (
		.in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_15_out));

	direct_interc direct_interc_16_ (
		.in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_16_out));

	direct_interc direct_interc_17_ (
		.in(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_17_out));

	direct_interc direct_interc_18_ (
		.in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_18_out));

	direct_interc direct_interc_19_ (
		.in(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_19_out));

	direct_interc direct_interc_20_ (
		.in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_20_out));

	direct_interc direct_interc_21_ (
		.in(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_21_out));

	direct_interc direct_interc_22_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_22_out));

	direct_interc direct_interc_23_ (
		.in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_23_out));

	direct_interc direct_interc_24_ (
		.in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_24_out));

	direct_interc direct_interc_25_ (
		.in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_25_out));

	direct_interc direct_interc_26_ (
		.in(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_26_out));

	direct_interc direct_interc_27_ (
		.in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_27_out));

	direct_interc direct_interc_28_ (
		.in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_28_out));

	direct_interc direct_interc_29_ (
		.in(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_29_out));

	direct_interc direct_interc_30_ (
		.in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_30_out));

	direct_interc direct_interc_31_ (
		.in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_31_out));

	direct_interc direct_interc_32_ (
		.in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_32_out));

	direct_interc direct_interc_33_ (
		.in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_33_out));

	direct_interc direct_interc_34_ (
		.in(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_34_out));

	direct_interc direct_interc_35_ (
		.in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_35_out));

	direct_interc direct_interc_36_ (
		.in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_36_out));

	direct_interc direct_interc_37_ (
		.in(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_37_out));

	direct_interc direct_interc_38_ (
		.in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_38_out));

	direct_interc direct_interc_39_ (
		.in(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_39_out));

	direct_interc direct_interc_40_ (
		.in(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_40_out));

	direct_interc direct_interc_41_ (
		.in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_41_out));

	direct_interc direct_interc_42_ (
		.in(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_42_out));

	direct_interc direct_interc_43_ (
		.in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_43_out));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
//`default_nettype none




